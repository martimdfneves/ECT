----------------------------------------------------------------------------------------------------------------------------------------------------------------
-- LSD.TOS, April 2018 (DO NOT REMOVE THIS LINE), VHDL 2008
--
-- Blop sound ROM (dual port, synchronous read). At 48kHz, this sound has a duration of about 85 miliseconds.
--
-- The blop sound was kindly put in the public domain by Mark DiAngelo (http://soundbible.com/2067-Blop.html).
--
-- Octave/matlab commands used to generate the data for the ROM:
--   x=wavread('Blop-Mark_DiAngelo-79054334.wav'); % read the .wav file
--   i=2496;                                       % index of the first sample we are interested in
--   y=round(65536*x(i:i+4095,1));                 % convert 4096 samples to integers (in this case, in the range -32767 to 32767)
--   y(end)=0;                                     % make sure the last sample is zero (silence)
--   save blop.txt y                               % save y
-- The 16-bit integers stored in the file blop.txt were then converted to hexadecimal and, after that, to VHDL.
--
-- A simple example of the use of the blop_sound_rom entity can be found in the file audio_example_tl.vhd
--

library IEEE;
use     IEEE.STD_LOGIC_1164.ALL;
use     IEEE.NUMERIC_STD.ALL;

entity blop_sound_rom is
  port
  (
    clock : in std_logic;

    addr0_0 : in  std_logic_vector(11 downto 0); -- sample number
    data0_1 : out std_logic_vector(15 downto 0); -- sample value (available with a delay of one clock cycle)

    addr1_0 : in  std_logic_vector(11 downto 0); -- sample number
    data1_1 : out std_logic_vector(15 downto 0)  -- sample value (available with a delay of one clock cycle)
  );
end blop_sound_rom;

architecture waveform_data of blop_sound_rom is
  --
  -- The sound samples (to be interpreted as 16-bit signed integers)
  --
  type rom_t is array(0 to 4095) of std_logic_vector(15 downto 0);
  constant WAVEFORM_DATA : rom_t :=
  (
    X"0004",X"0005",X"FFFE",X"FFFF",X"0009",X"0003",X"FFFC",X"FFF8",X"FFF7",X"FFF9",X"0001",X"0002",X"FFFF",X"FFFD",X"FFFE",X"FFF5",
    X"FFF2",X"FFF5",X"FFFD",X"FFF5",X"FFFE",X"FFFE",X"FFF8",X"FFF8",X"FFF6",X"FFEF",X"FFF7",X"FFFC",X"FFFE",X"FFFB",X"FFFA",X"FFF4",
    X"FFE8",X"FFE6",X"FFEB",X"FFF7",X"FFFD",X"0002",X"0003",X"FFF6",X"FFEF",X"FFE9",X"FFE8",X"FFEB",X"FFED",X"FFEC",X"FFE7",X"FFF0",
    X"FFF7",X"FFEF",X"FFE9",X"FFE1",X"FFDE",X"FFE7",X"FFE8",X"FFEA",X"FFE7",X"FFED",X"FFE9",X"FFEB",X"FFE5",X"FFDC",X"FFDE",X"FFDE",
    X"FFE2",X"FFD5",X"FFDA",X"FFD3",X"FFD7",X"FFD6",X"FFD7",X"FFCF",X"FFC1",X"FFBE",X"FFC3",X"FFCA",X"FFCE",X"FFCA",X"FFB7",X"FFB4",
    X"FFC0",X"FFD4",X"FFCE",X"FFCC",X"FFB9",X"FFB2",X"FFB4",X"FFB6",X"FFB5",X"FFC3",X"FFBF",X"FFB3",X"FFC1",X"FFC4",X"FFC9",X"FFCF",
    X"FFC2",X"FFAF",X"FF9F",X"FFAC",X"FFB6",X"FFAA",X"FFB2",X"FFBB",X"FFB9",X"FFB8",X"FFB0",X"FFAC",X"FFA0",X"FFB0",X"FFC6",X"FFBE",
    X"FFC1",X"FFB3",X"FF96",X"FF96",X"FFB6",X"FFC7",X"FFCB",X"FFC0",X"FFA3",X"FF7E",X"FF7E",X"FF8C",X"FFAB",X"FFC5",X"FFC4",X"FFC0",
    X"FFC2",X"FF97",X"FF91",X"FFA7",X"FFAC",X"FFCB",X"FFD8",X"FFC5",X"FFB6",X"FFC5",X"FFC5",X"FFC8",X"FFD4",X"FFD1",X"FFC5",X"FFB9",
    X"FFB3",X"FFC2",X"FFCC",X"FFD5",X"FFDB",X"FFD1",X"FFD9",X"FFCC",X"FFCE",X"FFD6",X"FFEB",X"FFFD",X"000D",X"FFF9",X"FFF3",X"FFD5",
    X"FFEA",X"FFF2",X"FFF4",X"001D",X"0003",X"0002",X"FFFC",X"0000",X"000C",X"0005",X"0012",X"0021",X"004C",X"0067",X"005C",X"003C",
    X"001A",X"0013",X"0025",X"0042",X"003C",X"0040",X"005B",X"001C",X"000A",X"0002",X"0017",X"0006",X"0002",X"0029",X"001E",X"FFB7",
    X"FF65",X"FF4E",X"FF26",X"FEE8",X"FE97",X"FE0A",X"FD2A",X"FC43",X"FB22",X"FA13",X"F8C2",X"F75C",X"F5BB",X"F40A",X"F275",X"F061",
    X"EE60",X"EC68",X"EA72",X"E832",X"E555",X"E0F9",X"DB79",X"D684",X"D398",X"D343",X"D46A",X"D45F",X"D2FF",X"D073",X"CDDE",X"CC0C",
    X"CB8C",X"CBF7",X"CC29",X"CC63",X"CCD1",X"CC87",X"CB95",X"CB34",X"CB2C",X"CAF1",X"CB93",X"CD24",X"CE6D",X"CE69",X"CDF0",X"CFA0",
    X"D1A8",X"D2F0",X"D4EC",X"D643",X"D7E2",X"D97E",X"DC02",X"DFDC",X"E074",X"E0E9",X"E3E7",X"E8E7",X"ECF1",X"EFC0",X"F231",X"F663",
    X"FA01",X"FEF1",X"0461",X"0934",X"0E34",X"13CC",X"1A29",X"1FF7",X"258B",X"29CA",X"2E63",X"33B8",X"38C1",X"3F1A",X"4466",X"48EF",
    X"4D4D",X"5219",X"56E1",X"5AF3",X"5F71",X"63AA",X"685B",X"6D93",X"70A6",X"736C",X"7588",X"766D",X"7795",X"7761",X"75B1",X"736C",
    X"704C",X"6C04",X"666C",X"5F81",X"57F0",X"4F63",X"4651",X"3C8B",X"3219",X"26E6",X"1B6E",X"102C",X"050D",X"F850",X"EBAE",X"E050",
    X"D471",X"C8BA",X"BDA7",X"B30A",X"A9A5",X"A258",X"9C23",X"9645",X"9286",X"9034",X"902B",X"922A",X"95D1",X"9A00",X"A02A",X"A7DA",
    X"B032",X"B995",X"C3E5",X"CE6D",X"DA00",X"E633",X"F28B",X"FF56",X"0C0C",X"18F6",X"25F4",X"32A2",X"3E28",X"4901",X"53AB",X"5D2D",
    X"65F7",X"6D2C",X"72A7",X"7601",X"7771",X"770E",X"750F",X"71AC",X"6C21",X"655C",X"5DCC",X"5482",X"4A12",X"3EB3",X"3268",X"25A4",
    X"18D2",X"0B13",X"FC79",X"EEB8",X"E1DD",X"D4E3",X"C861",X"BC6B",X"B16C",X"A851",X"A0D0",X"9A5C",X"95E9",X"936A",X"9296",X"9419",
    X"9739",X"9B06",X"A062",X"A790",X"B03F",X"B987",X"C367",X"CE23",X"D9CB",X"E611",X"F2AD",X"FF15",X"0B57",X"17AF",X"2410",X"3016",
    X"3B0A",X"454A",X"4EC6",X"56B9",X"5CF0",X"61D1",X"64D1",X"65E1",X"6580",X"638C",X"5FE8",X"5A74",X"5389",X"4B5C",X"425E",X"3884",
    X"2D6F",X"2160",X"14E8",X"086A",X"FC24",X"EFA5",X"E301",X"D6C1",X"CB25",X"C03E",X"B626",X"AD84",X"A6B4",X"A190",X"9E14",X"9C2E",
    X"9BD0",X"9D19",X"A016",X"A4B7",X"AADD",X"B21A",X"BA20",X"C396",X"CE5E",X"D975",X"E4C8",X"F090",X"FCB5",X"08BB",X"14D6",X"20D7",
    X"2C56",X"3748",X"41BC",X"4B2C",X"530B",X"5994",X"5ECB",X"6269",X"6449",X"6487",X"62F4",X"5FB7",X"5B11",X"553E",X"4DCF",X"44A9",
    X"3A8C",X"2FF2",X"2497",X"1874",X"0BFC",X"FF44",X"F28D",X"E621",X"D9D6",X"CDE7",X"C2CF",X"B8D4",X"B024",X"A8E7",X"A32D",X"9EFE",
    X"9C52",X"9B50",X"9C3C",X"9EC6",X"A2CD",X"A810",X"AEC2",X"B6F2",X"C018",X"C9CC",X"D41C",X"DF3F",X"EB0F",X"F73A",X"0327",X"0F0B",
    X"1AFC",X"267D",X"3154",X"3B51",X"4461",X"4C60",X"5324",X"585C",X"5BF5",X"5DFD",X"5E81",X"5D8B",X"5AFC",X"56EA",X"5139",X"4A10",
    X"41C3",X"3896",X"2E96",X"23C6",X"184C",X"0C5F",X"0048",X"F430",X"E846",X"DC84",X"D136",X"C688",X"BD11",X"B534",X"AED0",X"A981",
    X"A55B",X"A2C8",X"A232",X"A343",X"A5A3",X"A94E",X"AE64",X"B4D4",X"BC7D",X"C50D",X"CEA5",X"D8EA",X"E385",X"EE88",X"F9C2",X"053F",
    X"10EF",X"1C69",X"2749",X"3161",X"3ACB",X"4340",X"4A67",X"5055",X"551A",X"5863",X"59FF",X"5A45",X"5928",X"5649",X"51AC",X"4BD5",
    X"4503",X"3D12",X"33F7",X"29F0",X"1F5A",X"148D",X"0958",X"FDAC",X"F18B",X"E5AC",X"DA9D",X"D056",X"C6DF",X"BE44",X"B6A6",X"B053",
    X"AB5D",X"A7F0",X"A5D4",X"A542",X"A66F",X"A94E",X"AD9F",X"B2B7",X"B8BB",X"C004",X"C861",X"D190",X"DB41",X"E57D",X"F05D",X"FB61",
    X"0635",X"10E8",X"1B51",X"254A",X"2E9F",X"3707",X"3E59",X"44C8",X"4A4C",X"4E87",X"50FF",X"5203",X"51B0",X"4FDC",X"4CB7",X"486A",
    X"42FB",X"3C77",X"34E9",X"2C5F",X"2329",X"1952",X"0EFB",X"046E",X"F9D8",X"EF57",X"E531",X"DB8B",X"D29D",X"CAA7",X"C382",X"BD39",
    X"B830",X"B490",X"B276",X"B1BA",X"B23C",X"B40A",X"B6FF",X"BB2D",X"C049",X"C697",X"CE11",X"D653",X"DEF7",X"E7DA",X"F144",X"FB3A",
    X"051F",X"0EC3",X"1814",X"213C",X"2A00",X"31D6",X"38B3",X"3E83",X"430A",X"469F",X"4910",X"4A24",X"49DC",X"4859",X"45AB",X"419F",
    X"3C80",X"3671",X"2F91",X"27A7",X"1EDD",X"158C",X"0BD9",X"021E",X"F87B",X"EEEB",X"E550",X"DC0F",X"D391",X"CBF3",X"C547",X"BFA6",
    X"BB2F",X"B7E4",X"B5C3",X"B505",X"B59F",X"B77B",X"BA77",X"BE85",X"C38B",X"C95C",X"D025",X"D7DE",X"E03C",X"E8E3",X"F1E3",X"FB31",
    X"0482",X"0DCA",X"16E5",X"1FA0",X"27BB",X"2F1B",X"35C4",X"3B77",X"401B",X"439C",X"4604",X"470F",X"46CA",X"4587",X"4318",X"3F54",
    X"3A7A",X"34CC",X"2E3F",X"26BE",X"1EB7",X"162B",X"0D0E",X"039B",X"FA54",X"F14A",X"E885",X"DFE5",X"D7D9",X"D092",X"CA18",X"C49D",
    X"C067",X"BD49",X"BB47",X"BA77",X"BACC",X"BC4B",X"BEF9",X"C2BF",X"C780",X"CD07",X"D35B",X"DA65",X"E239",X"EA76",X"F314",X"FBDA",
    X"0480",X"0D1B",X"158A",X"1DB5",X"2548",X"2C27",X"3253",X"3792",X"3BC4",X"3EF8",X"412B",X"4226",X"41F2",X"408B",X"3E2C",X"3AC2",
    X"364B",X"30F1",X"2AAC",X"239C",X"1BEA",X"13D0",X"0B4B",X"029E",X"F9CD",X"F112",X"E890",X"E069",X"D8DB",X"D1F7",X"CBEF",X"C6CB",
    X"C2AD",X"BFAF",X"BDB9",X"BCD9",X"BD1C",X"BE89",X"C101",X"C453",X"C8A8",X"CDE0",X"D3D6",X"DA85",X"E1E4",X"E9AC",X"F1BB",X"FA05",
    X"025D",X"0AA6",X"12B6",X"1A7E",X"21D0",X"287A",X"2E77",X"339F",X"37F2",X"3B3B",X"3D6B",X"3EAC",X"3ED6",X"3DE0",X"3BF5",X"38FD",
    X"3506",X"302C",X"2A82",X"243B",X"1D49",X"15EC",X"0E1F",X"063E",X"FE2E",X"F62B",X"EE50",X"E6DB",X"DFBA",X"D958",X"D3B3",X"CED2",
    X"CAE2",X"C7D3",X"C5C9",X"C4CC",X"C4D0",X"C5D7",X"C7DC",X"CAB5",X"CE64",X"D2FF",X"D84B",X"DE27",X"E496",X"EB78",X"F292",X"F9DF",
    X"014C",X"08A4",X"0FC5",X"16A6",X"1D28",X"22FD",X"2827",X"2C9A",X"3050",X"332D",X"3508",X"360C",X"3629",X"3533",X"3343",X"309C",
    X"2D2B",X"28E8",X"23F8",X"1E62",X"183C",X"11BB",X"0AFB",X"0419",X"FD2E",X"F63F",X"EFA7",X"E95A",X"E380",X"DE1E",X"D99C",X"D5C8",
    X"D2B1",X"D07C",X"CF37",X"CEC9",X"CF39",X"D099",X"D2DB",X"D5C6",X"D971",X"DDCB",X"E2C6",X"E832",X"EE14",X"F454",X"FABF",X"013A",
    X"07A7",X"0E04",X"142C",X"19ED",X"1F46",X"240E",X"2822",X"2B88",X"2E2F",X"2FF4",X"30E6",X"30E6",X"301A",X"2E67",X"2BD9",X"2883",
    X"247A",X"1FDA",X"1A87",X"14B5",X"0E7D",X"0817",X"0179",X"FABF",X"F40D",X"ED8B",X"E756",X"E178",X"DC23",X"D77D",X"D381",X"D03B",
    X"CDCC",X"CC34",X"CB6D",X"CB9C",X"CC99",X"CE74",X"D122",X"D4A2",X"D8BE",X"DD6B",X"E2B7",X"E887",X"EE9D",X"F4FC",X"FB99",X"0233",
    X"08BB",X"0F21",X"1552",X"1B17",X"2053",X"2510",X"2929",X"2C85",X"2F1B",X"3103",X"320E",X"324F",X"31AE",X"3040",X"2DFE",X"2AFB",
    X"2745",X"22FD",X"1E11",X"18A8",X"12D5",X"0CB9",X"0660",X"0012",X"F9BB",X"F3A5",X"EDBA",X"E83B",X"E327",X"DEB0",X"DAD3",X"D7A1",
    X"D530",X"D378",X"D284",X"D260",X"D2F4",X"D442",X"D648",X"D90C",X"DC6B",X"E055",X"E4BC",X"E99D",X"EED7",X"F440",X"F9DD",X"FF8B",
    X"0533",X"0AA3",X"0FEB",X"14E4",X"1966",X"1D72",X"20E9",X"23C6",X"25F7",X"277F",X"2854",X"2875",X"27E6",X"2691",X"24AF",X"2211",
    X"1ED6",X"1B22",X"1709",X"126E",X"0DAD",X"08AD",X"0371",X"FE40",X"F91A",X"F427",X"EF6F",X"EB08",X"E713",X"E3A4",X"E0D0",X"DE89",
    X"DCED",X"DBF6",X"DB94",X"DBDC",X"DCD4",X"DE63",X"E094",X"E35C",X"E69E",X"EA4C",X"EE77",X"F2E0",X"F782",X"FC55",X"0135",X"0623",
    X"0AE7",X"0F72",X"13BC",X"17B8",X"1B46",X"1E42",X"20DA",X"22D2",X"2419",X"24CD",X"24FC",X"2473",X"2339",X"2174",X"1F1C",X"1C41",
    X"18E4",X"1513",X"10ED",X"0C7E",X"07D8",X"0317",X"FE30",X"F964",X"F4A9",X"F037",X"EBFE",X"E829",X"E4D7",X"E1EF",X"DF8D",X"DDC6",
    X"DC9C",X"DC04",X"DC16",X"DCBC",X"DDF3",X"DFBF",X"E211",X"E4D1",X"E810",X"EBB2",X"EFA5",X"F3E4",X"F852",X"FCD7",X"0162",X"05F2",
    X"0A55",X"0E89",X"1280",X"160C",X"1939",X"1BEC",X"1E21",X"1FD1",X"20FB",X"217B",X"2180",X"20EE",X"1FC1",X"1E18",X"1BE5",X"1935",
    X"1619",X"129D",X"0EC7",X"0AC7",X"0696",X"0242",X"FDEF",X"F9B2",X"F587",X"F199",X"EE06",X"EAAA",X"E7CF",X"E56D",X"E389",X"E237",
    X"E154",X"E0FB",X"E135",X"E215",X"E368",X"E526",X"E74B",X"E9EB",X"ECF9",X"F068",X"F40F",X"F7E7",X"FBE7",X"FFFE",X"03FC",X"07FC",
    X"0BC7",X"0F67",X"12B4",X"15A2",X"1833",X"1A52",X"1BF0",X"1D0B",X"1DA8",X"1DB5",X"1D3E",X"1C48",X"1ADA",X"18EF",X"168C",X"13C1",
    X"10B0",X"0D56",X"09B3",X"05E9",X"01FD",X"FDFF",X"FA0A",X"F638",X"F272",X"EEFD",X"EBE4",X"E914",X"E6B5",X"E4C3",X"E361",X"E261",
    X"E1F8",X"E20E",X"E2A9",X"E3B6",X"E545",X"E73B",X"E99B",X"EC61",X"EF69",X"F2CA",X"F658",X"FA01",X"FDC7",X"019F",X"0565",X"090B",
    X"0C8E",X"0FDB",X"12E9",X"1599",X"17DE",X"19BB",X"1B10",X"1BFE",X"1C70",X"1C60",X"1BD3",X"1AC6",X"1952",X"1779",X"1535",X"1296",
    X"0FB3",X"0C8E",X"0938",X"05BA",X"022E",X"FEA0",X"FB1D",X"F7C3",X"F491",X"F189",X"EEC9",X"EC5F",X"EA62",X"E8D1",X"E7B0",X"E701",
    X"E6D0",X"E703",X"E7A9",X"E8C6",X"EA43",X"EC29",X"EE6B",X"F0E6",X"F39C",X"F67E",X"F98E",X"FCD5",X"0019",X"0349",X"066D",X"0979",
    X"0C52",X"0EF4",X"114F",X"1357",X"14FD",X"164B",X"1724",X"1792",X"1796",X"1731",X"1646",X"14FD",X"1350",X"1156",X"0F0D",X"0C75",
    X"09A6",X"06B5",X"0395",X"007B",X"FD57",X"FA2B",X"F716",X"F442",X"F19B",X"EF47",X"ED32",X"EB6F",X"EA16",X"E91F",X"E894",X"E875",
    X"E8C6",X"E982",X"EA9A",X"EC15",X"EDE5",X"F013",X"F275",X"F50E",X"F7E2",X"FACD",X"FDCB",X"00E5",X"03E8",X"06E2",X"09BC",X"0C71",
    X"0EF9",X"1139",X"1328",X"14B9",X"15F5",X"16D6",X"1755",X"1769",X"1710",X"1651",X"1537",X"13AF",X"11EE",X"0FC5",X"0D68",X"0ADE",
    X"0815",X"053A",X"0233",X"FF32",X"FC3C",X"F942",X"F677",X"F3DB",X"F17A",X"EF4B",X"ED8B",X"EC07",X"EAED",X"EA2C",X"E9C5",X"E9D7",
    X"EA3E",X"EB0A",X"EC30",X"EDAF",X"EF7D",X"F189",X"F3D4",X"F65A",X"F906",X"FBCE",X"FEAE",X"0184",X"045C",X"0720",X"09BF",X"0C30",
    X"0E6C",X"1066",X"121D",X"1379",X"1484",X"1530",X"1571",X"155B",X"14FD",X"142E",X"130F",X"1197",X"0FD2",X"0DDA",X"0BB9",X"094A",
    X"06C5",X"0422",X"0188",X"FEDA",X"FC47",X"F9BB",X"F757",X"F529",X"F32F",X"F185",X"F029",X"EF11",X"EE4E",X"EDDC",X"EDC1",X"EE06",
    X"EEAC",X"EFA5",X"F0F1",X"F275",X"F439",X"F634",X"F86D",X"FAB8",X"FD2A",X"FF97",X"0225",X"049B",X"06FD",X"0938",X"0B57",X"0D44",
    X"0EF2",X"105B",X"117A",X"123B",X"12C6",X"12FB",X"12DA",X"126E",X"11B0",X"1097",X"0F33",X"0D8B",X"0BAE",X"09A2",X"0766",X"051B",
    X"02B2",X"003F",X"FDBB",X"FB58",X"F90A",X"F6DA",X"F4DB",X"F311",X"F183",X"F03E",X"EF40",X"EE82",X"EE2A",X"EE26",X"EE6B",X"EEF2",
    X"EFD4",X"F101",X"F263",X"F411",X"F5E3",X"F7D9",X"F9FC",X"FC38",X"FE7A",X"00D9",X"0325",X"0565",X"0785",X"097E",X"0B47",X"0CE1",
    X"0E4C",X"0F6D",X"1047",X"10D2",X"1107",X"10EF",X"108A",X"0FE0",X"0EFB",X"0DC3",X"0C5B",X"0AB5",X"08DC",X"06D7",X"04B8",X"0288",
    X"003D",X"FE05",X"FBDC",X"F9BB",X"F7B1",X"F5CF",X"F421",X"F2C1",X"F180",X"F097",X"EFE6",X"EF7F",X"EF6D",X"EF9A",X"F020",X"F0EF",
    X"F1F3",X"F341",X"F4C0",X"F66C",X"F850",X"FA44",X"FC6B",X"FE9E",X"00D5",X"02F8",X"0502",X"06EF",X"08D8",X"0A91",X"0C13",X"0D58",
    X"0E60",X"0F35",X"0FB5",X"0FDD",X"0FC5",X"0F6D",X"0ED9",X"0DF3",X"0CCB",X"0B76",X"09DC",X"0817",X"062E",X"0419",X"01F6",X"FFCF",
    X"FDB7",X"FB9D",X"F98E",X"F7A6",X"F5D6",X"F439",X"F2D7",X"F1B2",X"F0DD",X"F03B",X"EFDD",X"EFC2",X"F003",X"F07F",X"F142",X"F23F",
    X"F37F",X"F4DF",X"F687",X"F859",X"FA42",X"FC41",X"FE5B",X"0077",X"0295",X"04A2",X"06A1",X"088C",X"0A4E",X"0BC4",X"0D0E",X"0E26",
    X"0EFF",X"0F96",X"0FEF",X"0FEF",X"0FC2",X"0F47",X"0E84",X"0D94",X"0C5F",X"0AFB",X"096C",X"07BD",X"05DE",X"03F1",X"01FF",X"FFF7",
    X"FDF8",X"FC0B",X"FA32",X"F864",X"F6D1",X"F568",X"F435",X"F338",X"F267",X"F209",X"F1CA",X"F1D3",X"F214",X"F2A8",X"F36D",X"F46F",
    X"F5A4",X"F70D",X"F8AC",X"FA61",X"FC38",X"FE17",X"000B",X"01F6",X"03D8",X"05AA",X"076F",X"0919",X"0A8B",X"0BD4",X"0CF5",X"0DD1",
    X"0E80",X"0EE0",X"0F04",X"0EE5",X"0E7D",X"0DE3",X"0D09",X"0BFA",X"0AB5",X"0946",X"07B4",X"05F0",X"0434",X"0252",X"0060",X"FE81",
    X"FCAA",X"FAE5",X"F935",X"F7A1",X"F634",X"F503",X"F401",X"F33E",X"F2C5",X"F277",X"F279",X"F2AA",X"F323",X"F3D7",X"F4B7",X"F5D4",
    X"F714",X"F884",X"FA0E",X"FBB8",X"FD78",X"FF3B",X"0106",X"02D4",X"0496",X"064C",X"07D4",X"093D",X"0A94",X"0BBE",X"0CA9",X"0D5A",
    X"0DDA",X"0E07",X"0E14",X"0DD5",X"0D61",X"0CB4",X"0BC7",X"0A9D",X"0943",X"07CD",X"0633",X"0487",X"02C2",X"00EE",X"FF2B",X"FD60",
    X"FB9B",X"F9E4",X"F855",X"F6EE",X"F5B2",X"F49C",X"F3B1",X"F30F",X"F29F",X"F272",X"F279",X"F2B6",X"F338",X"F3E6",X"F4D2",X"F5F1",
    X"F736",X"F893",X"FA13",X"FBBC",X"FD6F",X"FF30",X"00F4",X"02AE",X"0451",X"05E2",X"075B",X"08BD",X"09EB",X"0AEB",X"0BBE",X"0C64",
    X"0CD4",X"0D07",X"0D00",X"0CBB",X"0C37",X"0B91",X"0AB7",X"099F",X"0868",X"06FA",X"0589",X"03F1",X"023E",X"008D",X"FEDD",X"FD28",
    X"FB7E",X"F9EA",X"F86D",X"F724",X"F5F7",X"F4F1",X"F421",X"F37D",X"F311",X"F2D9",X"F302",X"F338",X"F3C0",X"F46D",X"F54B",X"F656",
    X"F780",X"F8C7",X"FA32",X"FBC1",X"FD5B",X"FEFE",X"00A1",X"0240",X"03D8",X"0567",X"06C7",X"0815",X"093A",X"0A41",X"0B08",X"0BA7",
    X"0C0C",X"0C42",X"0C40",X"0C01",X"0BAA",X"0B13",X"0A50",X"095E",X"0844",X"0718",X"05CA",X"0453",X"02CF",X"0157",X"FFE5",X"FE64",
    X"FCE7",X"FB7E",X"FA2B",X"F8F6",X"F7E0",X"F6EC",X"F62B",X"F595",X"F539",X"F517",X"F513",X"F549",X"F5A7",X"F632",X"F6F0",X"F7DC",
    X"F8D9",X"F9FE",X"FB3D",X"FC7D",X"FDDF",X"FF53",X"00BC",X"0230",X"038A",X"04DC",X"0623",X"073E",X"0842",X"092B",X"09DA",X"0A70",
    X"0AD5",X"0B04",X"0B1A",X"0AFF",X"0AAA",X"0A4A",X"09AF",X"08EA",X"0805",X"0708",X"05F6",X"04D1",X"0395",X"0250",X"010D",X"FFC8",
    X"FE95",X"FD60",X"FC45",X"FB2D",X"FA4D",X"F978",X"F8C9",X"F849",X"F7E7",X"F7BE",X"F7BA",X"F7BC",X"F804",X"F862",X"F8E8",X"F98E",
    X"FA48",X"FB26",X"FC16",X"FD23",X"FE2C",X"FF4D",X"0069",X"0182",X"0297",X"039B",X"0489",X"0569",X"062A",X"06C9",X"0754",X"07BD",
    X"0801",X"0827",X"0822",X"0801",X"07AE",X"073E",X"06AA",X"060D",X"0551",X"0479",X"0395",X"0297",X"019F",X"009F",X"FF9B",X"FE8E",
    X"FD9C",X"FCBC",X"FBDC",X"FB22",X"FA80",X"F9F3",X"F97A",X"F932",X"F90C",X"F91A",X"F932",X"F962",X"F9A7",X"FA20",X"FA9E",X"FB3F",
    X"FBFB",X"FCC3",X"FD95",X"FE76",X"FF58",X"0048",X"012F",X"0218",X"02F3",X"03C8",X"046E",X"0524",X"05B3",X"0623",X"067F",X"06BC",
    X"06DF",X"06E4",X"06C0",X"0681",X"062C",X"05BC",X"0531",X"049F",X"03F3",X"0340",X"026F",X"019C",X"00BA",X"FFDE",X"FEFA",X"FE20",
    X"FD50",X"FC79",X"FBC1",X"FB17",X"FA8C",X"FA19",X"F9B9",X"F978",X"F95D",X"F954",X"F96A",X"F97A",X"F9BB",X"FA19",X"FA8C",X"FAFE",
    X"FB8D",X"FC28",X"FCCC",X"FD7D",X"FE35",X"FEEA",X"FFA4",X"0063",X"0111",X"01B1",X"0237",X"02B9",X"0329",X"0395",X"03D8",X"0409",
    X"042D",X"0438",X"0432",X"0417",X"03E5",X"03B0",X"0363",X"030E",X"02B7",X"024B",X"01D9",X"015E",X"00E0",X"006C",X"FFFE",X"FF8E",
    X"FF2D",X"FED8",X"FE87",X"FE3D",X"FE0C",X"FDDF",X"FDBB",X"FDC2",X"FDCB",X"FDF6",X"FE2C",X"FE66",X"FEB0",X"FF12",X"FF75",X"FFE3",
    X"0043",X"00B8",X"0126",X"018F",X"01F8",X"024B",X"0297",X"02E6",X"0322",X"0349",X"0366",X"036F",X"0366",X"0351",X"033D",X"0303",
    X"02D2",X"027A",X"021C",X"01AE",X"0138",X"00B8",X"002F",X"FFB4",X"FF2D",X"FEB4",X"FE40",X"FDD2",X"FD6D",X"FD11",X"FCB7",X"FC82",
    X"FC50",X"FC38",X"FC31",X"FC33",X"FC4A",X"FC7B",X"FCBA",X"FD11",X"FD7F",X"FDFA",X"FE73",X"FEFA",X"FF8E",X"0026",X"00BC",X"0159",
    X"01EF",X"0281",X"030A",X"0387",X"0400",X"0458",X"04B4",X"04EE",X"0524",X"053C",X"053F",X"0524",X"04FB",X"04B6",X"0480",X"0412",
    X"0399",X"030E",X"0286",X"01F8",X"0147",X"009F",X"FFF9",X"FF56",X"FEC6",X"FE1A",X"FD8A",X"FD13",X"FC91",X"FC31",X"FBE3",X"FBA6",
    X"FB80",X"FB75",X"FB75",X"FB96",X"FBCE",X"FC0D",X"FC62",X"FCD0",X"FD50",X"FDE4",X"FE7C",X"FF20",X"FFD8",X"0082",X"0126",X"01CE",
    X"026B",X"0305",X"0397",X"0419",X"0485",X"04CA",X"0516",X"0538",X"0551",X"054C",X"052D",X"04EE",X"049B",X"0438",X"03C6",X"033D",
    X"02A3",X"0208",X"0157",X"0098",X"FFDC",X"FF19",X"FE68",X"FDB0",X"FCFD",X"FC59",X"FBCC",X"FB46",X"FAD6",X"FA73",X"FA27",X"FA01",
    X"F9DB",X"F9E4",X"FA05",X"FA34",X"FA7C",X"FAE1",X"FB65",X"FBE0",X"FC79",X"FD31",X"FDFA",X"FEAB",X"FF5F",X"001B",X"00D7",X"019A",
    X"0252",X"02FF",X"0395",X"041D",X"049F",X"0504",X"0560",X"059A",X"05D3",X"05E2",X"05CE",X"05A8",X"056E",X"0524",X"04BF",X"0444",
    X"03B6",X"0320",X"0278",X"01C9",X"011D",X"005E",X"FFA4",X"FEF5",X"FE58",X"FDB3",X"FD1C",X"FC94",X"FC21",X"FBC5",X"FB67",X"FB3D",
    X"FB12",X"FB07",X"FB12",X"FB2F",X"FB6A",X"FBA8",X"FC06",X"FC76",X"FCF2",X"FD8A",X"FE13",X"FE99",X"FF32",X"FFC6",X"005E",X"00EB",
    X"0172",X"01F8",X"0262",X"02C9",X"0329",X"0366",X"039E",X"03C6",X"03D6",X"03DA",X"03CD",X"03A4",X"037E",X"0334",X"02D4",X"0278",
    X"0208",X"019A",X"011F",X"0096",X"0024",X"FFA2",X"FF27",X"FEB0",X"FE3B",X"FDDB",X"FD88",X"FD40",X"FD06",X"FCDB",X"FCC0",X"FCB7",
    X"FCBC",X"FCD5",X"FCFF",X"FD35",X"FD78",X"FDD2",X"FE2C",X"FE8C",X"FF0C",X"FF8B",X"0009",X"007B",X"00F2",X"016B",X"01D9",X"024B",
    X"02A3",X"02E4",X"032E",X"0358",X"0373",X"0387",X"0387",X"037C",X"0363",X"0329",X"02E8",X"0295",X"0242",X"01DD",X"0176",X"0102",
    X"0082",X"0009",X"FF90",X"FF19",X"FEAB",X"FE35",X"FDC9",X"FD66",X"FD18",X"FCDE",X"FC9F",X"FC79",X"FC69",X"FC5E",X"FC7B",X"FC86",
    X"FCBA",X"FCED",X"FD31",X"FD88",X"FDEF",X"FE5D",X"FEBF",X"FF27",X"FFB4",X"0031",X"00A1",X"011D",X"0179",X"01D2",X"022C",X"026B",
    X"02A7",X"02D6",X"0305",X"030E",X"0310",X"0301",X"02E1",X"02B2",X"0278",X"0235",X"01E9",X"0182",X"011D",X"00B6",X"004C",X"FFE3",
    X"FF68",X"FF05",X"FEA9",X"FE42",X"FDF4",X"FDA5",X"FD57",X"FD25",X"FCF4",X"FCDB",X"FCCE",X"FCCE",X"FCE9",X"FD0F",X"FD45",X"FD88",
    X"FDD9",X"FE32",X"FE8E",X"FEF3",X"FF6E",X"FFE7",X"0067",X"00E5",X"0164",X"01D7",X"0254",X"02B7",X"0310",X"035F",X"0395",X"03CF",
    X"03FC",X"0405",X"0409",X"0403",X"03DF",X"03A7",X"0363",X"0313",X"02BB",X"024B",X"01D0",X"0162",X"00D3",X"0045",X"FFBD",X"FF41",
    X"FEB2",X"FE30",X"FDAE",X"FD3C",X"FCDE",X"FC79",X"FC33",X"FBF0",X"FBC5",X"FBAD",X"FBA4",X"FBAF",X"FBC8",X"FBF7",X"FC38",X"FC82",
    X"FCD7",X"FD3E",X"FDB3",X"FE2E",X"FEB0",X"FF2B",X"FFBD",X"0045",X"00E2",X"016D",X"01FD",X"026D",X"02DF",X"0340",X"038E",X"03D3",
    X"0409",X"0419",X"0426",X"0419",X"0410",X"03E1",X"03AB",X"036C",X"0322",X"02D6",X"025F",X"01F6",X"017F",X"0100",X"0084",X"0000",
    X"FF82",X"FF05",X"FE90",X"FE20",X"FDB7",X"FD64",X"FD16",X"FCDE",X"FC9F",X"FC7D",X"FC74",X"FC67",X"FC7D",X"FC98",X"FCBE",X"FCFB",
    X"FD47",X"FD9E",X"FDFF",X"FE6A",X"FED4",X"FF51",X"FFC1",X"002B",X"00A1",X"0114",X"016D",X"01C9",X"0213",X"025D",X"0297",X"02BB",
    X"02CF",X"02ED",X"02EA",X"02DF",X"02C0",X"0293",X"0256",X"0208",X"01B3",X"0160",X"00F2",X"0080",X"0019",X"FFAD",X"FF36",X"FEBF",
    X"FE4B",X"FDE4",X"FD8F",X"FD35",X"FCE9",X"FCB3",X"FC7F",X"FC5E",X"FC47",X"FC45",X"FC55",X"FC70",X"FCA6",X"FCE2",X"FD1C",X"FD6D",
    X"FDC2",X"FE27",X"FE8C",X"FF00",X"FF77",X"FFEE",X"0063",X"00E0",X"0160",X"01C3",X"0225",X"027F",X"02DD",X"031C",X"0346",X"0373",
    X"037C",X"0387",X"0381",X"0371",X"0349",X"0327",X"02E6",X"02A7",X"0262",X"0208",X"01A5",X"0145",X"00DE",X"0069",X"0007",X"FF99",
    X"FF30",X"FECF",X"FE7A",X"FE29",X"FDDB",X"FDAE",X"FD7A",X"FD62",X"FD52",X"FD57",X"FD6D",X"FD8F",X"FDA7",X"FDDF",X"FE20",X"FE52",
    X"FE99",X"FEF3",X"FF46",X"FFB2",X"0009",X"0069",X"00D0",X"011D",X"0174",X"01D0",X"020F",X"024B",X"028A",X"02AC",X"02C7",X"02CD",
    X"02D2",X"02BE",X"02B0",X"027A",X"0242",X"0201",X"01BE",X"0164",X"0116",X"00BF",X"0067",X"FFFC",X"FF9D",X"FF39",X"FEDA",X"FE81",
    X"FE2C",X"FDDD",X"FD9C",X"FD66",X"FD45",X"FD2C",X"FD28",X"FD28",X"FD31",X"FD47",X"FD6F",X"FD9E",X"FDE4",X"FE23",X"FE64",X"FEBB",
    X"FF12",X"FF68",X"FFD3",X"0024",X"0084",X"00D3",X"0118",X"016B",X"01B7",X"01E4",X"021A",X"023E",X"0252",X"025F",X"025F",X"0256",
    X"0237",X"0211",X"01DB",X"019A",X"0149",X"0100",X"00AA",X"0048",X"FFE5",X"FF7E",X"FF1E",X"FEC4",X"FE61",X"FE0C",X"FDB3",X"FD64",
    X"FD1F",X"FCF0",X"FCCC",X"FCB1",X"FCA3",X"FCAA",X"FCAF",X"FCC5",X"FCF6",X"FD28",X"FD62",X"FDB7",X"FE11",X"FE76",X"FEE3",X"FF48",
    X"FFB4",X"0024",X"0092",X"00FB",X"0160",X"01C5",X"021A",X"0281",X"02C0",X"02F1",X"0329",X"0342",X"0349",X"034D",X"0337",X"030A",
    X"02CB",X"027D",X"0237",X"01E6",X"0176",X"00FD",X"008B",X"0010",X"FF8E",X"FF07",X"FE87",X"FE0A",X"FD9E",X"FD2C",X"FCC5",X"FC70",
    X"FC12",X"FBCC",X"FBA8",X"FB80",X"FB77",X"FB79",X"FB99",X"FBBA",X"FBF7",X"FC4C",X"FC9F",X"FCF8",X"FD74",X"FDF6",X"FE87",X"FF22",
    X"FFB6",X"004A",X"00E0",X"0176",X"0206",X"0288",X"030C",X"037E",X"03EE",X"044D",X"0485",X"04A6",X"04C6",X"04CA",X"04BA",X"0492",
    X"0463",X"0410",X"03B0",X"034D",X"02D8",X"0259",X"01C5",X"0131",X"0094",X"000B",X"FF68",X"FED8",X"FE4F",X"FDD9",X"FD59",X"FCE0",
    X"FC70",X"FC1B",X"FBD1",X"FBA4",X"FB75",X"FB70",X"FB79",X"FB87",X"FBB1",X"FBF7",X"FC43",X"FC9D",X"FCF8",X"FD78",X"FDF4",X"FE81",
    X"FF0C",X"FFA6",X"0036",X"00BC",X"014E",X"01CE",X"0247",X"02B2",X"0322",X"036F",X"03BD",X"03F7",X"0412",X"0429",X"0424",X"0419",
    X"0403",X"03D1",X"038C",X"0337",X"02CF",X"0266",X"01F4",X"017F",X"00F9",X"0075",X"FFE7",X"FF65",X"FEE1",X"FE64",X"FDF1",X"FD8A",
    X"FD2C",X"FCD7",X"FC9D",X"FC55",X"FC3A",X"FC2D",X"FC35",X"FC3C",X"FC60",X"FC9F",X"FCE9",X"FD3C",X"FDAA",X"FE15",X"FE8E",X"FF03",
    X"FF82",X"0007",X"008B",X"010B",X"0176",X"01E9",X"023E",X"02A7",X"0303",X"0349",X"038E",X"03B0",X"03B6",X"03BB",X"039E",X"037C",
    X"034B",X"0301",X"02B5",X"0247",X"01D2",X"0157",X"00E7",X"005C",X"FFD5",X"FF4D",X"FEB9",X"FE37",X"FDC0",X"FD50",X"FCEB",X"FC86",
    X"FC47",X"FC00",X"FBCE",X"FBA8",X"FBB1",X"FBB1",X"FBCA",X"FBF7",X"FC2D",X"FC74",X"FCE2",X"FD47",X"FDC4",X"FE56",X"FED6",X"FF61",
    X"FFF7",X"008F",X"0123",X"01B5",X"023E",X"02B7",X"0325",X"0399",X"03F3",X"0434",X"046A",X"0485",X"049D",X"04AB",X"049B",X"0479",
    X"043D",X"03F3",X"0392",X"0329",X"02B2",X"0237",X"01BA",X"0116",X"0084",X"FFE7",X"FF4F",X"FEC2",X"FE2E",X"FDB0",X"FD31",X"FCC9",
    X"FC62",X"FC0F",X"FBBA",X"FB96",X"FB75",X"FB6C",X"FB7B",X"FB99",X"FBCE",X"FC0B",X"FC5E",X"FCCC",X"FD39",X"FDC0",X"FE4B",X"FEE6",
    X"FF7A",X"001F",X"00CE",X"015E",X"01F8",X"0286",X"0305",X"038A",X"03F5",X"0453",X"04A4",X"04E0",X"0518",X"052A",X"0524",X"0509",
    X"04E7",X"04A8",X"045C",X"0405",X"0381",X"0303",X"0288",X"01F2",X"015B",X"00B1",X"000B",X"FF58",X"FEC6",X"FE27",X"FD86",X"FD04",
    X"FC76",X"FC06",X"FBA6",X"FB53",X"FB20",X"FB02",X"FAEC",X"FAEA",X"FB02",X"FB31",X"FB72",X"FBBC",X"FC1F",X"FC9A",X"FD0F",X"FD91",
    X"FE15",X"FEB0",X"FF48",X"FFE1",X"0077",X"011D",X"01A3",X"022A",X"02B9",X"0330",X"03A2",X"03EC",X"043F",X"0470",X"0499",X"04B4",
    X"04BD",X"04AD",X"0489",X"045A",X"0419",X"03CB",X"036C",X"0310",X"02A5",X"0223",X"01B3",X"011D",X"0094",X"0000",X"FF73",X"FEFC",
    X"FE76",X"FE03",X"FD95",X"FD28",X"FCC9",X"FC86",X"FC55",X"FC31",X"FC18",X"FC0B",X"FC16",X"FC28",X"FC47",X"FC84",X"FCC9",X"FD13",
    X"FD54",X"FDAC",X"FE1A",X"FE83",X"FEF3",X"FF56",X"FFC8",X"0026",X"0096",X"00F7",X"015E",X"01AA",X"01FF",X"023E",X"0271",X"0297",
    X"02B2",X"02BE",X"02B9",X"02A5",X"028A",X"0268",X"0223",X"01F2",X"019C",X"015B",X"010F",X"00BF",X"006C",X"000D",X"FFB8",X"FF5F",
    X"FF12",X"FEBD",X"FE71",X"FE32",X"FDFC",X"FDC2",X"FDA5",X"FD8A",X"FD76",X"FD76",X"FD7A",X"FD93",X"FDAC",X"FDE4",X"FE11",X"FE3B",
    X"FE87",X"FECD",X"FF1E",X"FF6A",X"FFBB",X"0010",X"005E",X"00A4",X"0104",X"0143",X"0198",X"01D2",X"0206",X"022C",X"0256",X"0266",
    X"0283",X"0288",X"028A",X"028C",X"026D",X"0249",X"0215",X"01E0",X"019F",X"0155",X"0114",X"00C5",X"0072",X"001B",X"FFD1",X"FF7E",
    X"FF29",X"FEEF",X"FEA9",X"FE6F",X"FE3B",X"FE15",X"FE08",X"FDE6",X"FDDD",X"FDE2",X"FDF6",X"FDFA",X"FE1E",X"FE3D",X"FE5F",X"FE8A",
    X"FEBD",X"FEFA",X"FF34",X"FF73",X"FFCA",X"0014",X"005A",X"00AD",X"0106",X"015B",X"01A5",X"01CE",X"0208",X"0230",X"0259",X"0274",
    X"0281",X"0283",X"027D",X"0268",X"024B",X"022C",X"01FD",X"01D4",X"019F",X"0164",X"0126",X"00E2",X"0092",X"0045",X"FFFC",X"FFAD",
    X"FF5F",X"FF03",X"FEB4",X"FE71",X"FE35",X"FE08",X"FDCB",X"FDA7",X"FD8A",X"FD7A",X"FD7D",X"FD7A",X"FD7F",X"FD9C",X"FDBE",X"FDD6",
    X"FDF6",X"FE1C",X"FE58",X"FE8A",X"FEBD",X"FF00",X"FF3B",X"FF7C",X"FFC6",X"0009",X"004C",X"0086",X"00C7",X"00F7",X"012F",X"0152",
    X"0169",X"017F",X"0193",X"01A8",X"01AA",X"01A8",X"01A8",X"019A",X"0179",X"0170",X"0155",X"0135",X"0114",X"00F9",X"00D0",X"009F",
    X"0077",X"004C",X"0014",X"FFF7",X"FFC3",X"FF9D",X"FF85",X"FF71",X"FF51",X"FF3B",X"FF22",X"FF15",X"FF12",X"FF05",X"FF17",X"FF1B",
    X"FF29",X"FF30",X"FF46",X"FF5F",X"FF7A",X"FF90",X"FFA6",X"FFC8",X"FFF5",X"0012",X"0036",X"004C",X"0069",X"0086",X"0092",X"00A6",
    X"00C1",X"00B3",X"00A1",X"00A6",X"009B",X"0096",X"0089",X"0080",X"0063",X"0055",X"0043",X"002D",X"002B",X"0024",X"001B",X"FFFE",
    X"FFEE",X"FFCF",X"FFD3",X"FFBF",X"FFAD",X"FFA9",X"FF99",X"FF97",X"FF8E",X"FF90",X"FF99",X"FF92",X"FF99",X"FFA9",X"FFBB",X"FFC3",
    X"FFD8",X"FFE5",X"000B",X"001F",X"003A",X"0057",X"0063",X"006E",X"0098",X"00A4",X"00BA",X"00C5",X"00C7",X"00E5",X"00F2",X"00F9",
    X"00FD",X"00FD",X"010D",X"0102",X"0102",X"0100",X"00F0",X"00D5",X"00C1",X"00A6",X"0092",X"0089",X"0065",X"0055",X"002D",X"001B",
    X"0000",X"FFEE",X"FFCF",X"FFBF",X"FFA9",X"FF94",X"FF85",X"FF73",X"FF68",X"FF51",X"FF5A",X"FF5A",X"FF5C",X"FF5F",X"FF5F",X"FF68",
    X"FF73",X"FF90",X"FFA2",X"FFB8",X"FFD1",X"FFEC",X"0004",X"001D",X"003F",X"005C",X"007B",X"00A1",X"00B3",X"00D7",X"00EB",X"0108",
    X"0114",X"012F",X"0150",X"0157",X"0164",X"016D",X"0170",X"0174",X"016D",X"016B",X"0150",X"0149",X"0145",X"0133",X"0123",X"010B",
    X"00F9",X"00D9",X"00B6",X"0098",X"0080",X"005E",X"0041",X"0028",X"0007",X"FFF5",X"FFD8",X"FFC3",X"FFA6",X"FF9D",X"FF97",X"FF92",
    X"FF99",X"FF9B",X"FF95",X"FF9B",X"FFA0",X"FFB0",X"FFB2",X"FFBE",X"FFD8",X"FFF1",X"000D",X"000F",X"001A",X"0032",X"004E",X"0056",
    X"005D",X"006A",X"0079",X"0077",X"0080",X"0086",X"008E",X"0082",X"0077",X"006F",X"0061",X"004A",X"0040",X"0024",X"0014",X"FFF0",
    X"FFD2",X"FFB5",X"FF93",X"FF81",X"FF62",X"FF4F",X"FF2E",X"FF13",X"FEF0",X"FED5",X"FEBE",X"FEB4",X"FE98",X"FE93",X"FE95",X"FE8F",
    X"FE93",X"FE92",X"FE98",X"FEB0",X"FEC2",X"FED2",X"FEED",X"FF0A",X"FF1E",X"FF43",X"FF6B",X"FF8E",X"FFC0",X"FFE9",X"0017",X"0041",
    X"0077",X"00A5",X"00DB",X"010E",X"0138",X"0156",X"017C",X"019F",X"01C3",X"01C9",X"01D5",X"01EC",X"01F8",X"01F0",X"01E4",X"01DC",
    X"01CC",X"01BB",X"019A",X"0187",X"0163",X"0136",X"0111",X"00E2",X"00AF",X"0071",X"003A",X"0010",X"FFDE",X"FFA5",X"FF77",X"FF4E",
    X"FF1C",X"FEFF",X"FEDF",X"FEC1",X"FEAA",X"FE99",X"FE84",X"FE7A",X"FE72",X"FE76",X"FE79",X"FE7F",X"FE7C",X"FE99",X"FEA7",X"FEB7",
    X"FED4",X"FEFC",X"FF19",X"FF3F",X"FF71",X"FFA4",X"FFC4",X"FFEE",X"001B",X"0042",X"0071",X"0092",X"00B7",X"00D0",X"00F3",X"0109",
    X"0121",X"0127",X"0136",X"013B",X"0142",X"013D",X"0138",X"0134",X"011B",X"00FF",X"00E9",X"00D3",X"00B3",X"0090",X"0077",X"0056",
    X"0035",X"0015",X"FFF6",X"FFD9",X"FFB9",X"FF9D",X"FF80",X"FF6C",X"FF4F",X"FF44",X"FF33",X"FF26",X"FF23",X"FF24",X"FF26",X"FF2D",
    X"FF36",X"FF44",X"FF4D",X"FF5A",X"FF74",X"FF88",X"FFA3",X"FFBD",X"FFDB",X"FFF5",X"0012",X"0031",X"0048",X"0062",X"0070",X"0081",
    X"009D",X"00A8",X"00B8",X"00C2",X"00C8",X"00C5",X"00CB",X"00C7",X"00BF",X"00B9",X"00B4",X"00A3",X"0094",X"007D",X"0066",X"004C",
    X"0038",X"001F",X"0007",X"FFF3",X"FFD9",X"FFC4",X"FFAB",X"FF97",X"FF8A",X"FF76",X"FF76",X"FF65",X"FF5B",X"FF58",X"FF55",X"FF52",
    X"FF56",X"FF5D",X"FF65",X"FF72",X"FF81",X"FF92",X"FFA6",X"FFBD",X"FFD5",X"FFE7",X"0005",X"001C",X"0034",X"0048",X"005E",X"0076",
    X"0088",X"0098",X"00AD",X"00B6",X"00C1",X"00C6",X"00C6",X"00C9",X"00C3",X"00BB",X"00AF",X"009E",X"0092",X"007B",X"006A",X"0057",
    X"0043",X"0029",X"0013",X"FFFE",X"FFEB",X"FFD1",X"FFB8",X"FFA6",X"FF8D",X"FF7D",X"FF6D",X"FF60",X"FF55",X"FF50",X"FF4B",X"FF4A",
    X"FF48",X"FF4F",X"FF51",X"FF5A",X"FF67",X"FF78",X"FF86",X"FF99",X"FFAD",X"FFC5",X"FFDA",X"FFF5",X"000D",X"0022",X"0036",X"004D",
    X"0062",X"0073",X"0081",X"0092",X"00A0",X"00A7",X"00B4",X"00BC",X"00BE",X"00B9",X"00B5",X"00B5",X"00AB",X"00A2",X"0094",X"0088",
    X"0078",X"0064",X"004F",X"003F",X"002A",X"0014",X"FFFE",X"FFED",X"FFD5",X"FFBD",X"FFAE",X"FF9B",X"FF88",X"FF7C",X"FF71",X"FF66",
    X"FF5F",X"FF5C",X"FF59",X"FF5A",X"FF5E",X"FF68",X"FF6E",X"FF7A",X"FF87",X"FF95",X"FFA7",X"FFB7",X"FFC7",X"FFDD",X"FFEF",X"0001",
    X"0014",X"0027",X"0038",X"0045",X"0057",X"0063",X"006E",X"0078",X"0081",X"0084",X"0089",X"008D",X"008E",X"0088",X"0085",X"0080",
    X"0075",X"0068",X"005C",X"004D",X"0043",X"0031",X"001E",X"0015",X"0002",X"FFF4",X"FFE9",X"FFD9",X"FFCD",X"FFC0",X"FFBA",X"FFB4",
    X"FFAD",X"FFAB",X"FFA5",X"FFA6",X"FFA7",X"FFAA",X"FFAA",X"FFB2",X"FFB7",X"FFC1",X"FFC9",X"FFD6",X"FFE0",X"FFEB",X"FFF8",X"0005",
    X"0014",X"0020",X"002C",X"0036",X"0043",X"004A",X"0053",X"005B",X"0061",X"0065",X"0068",X"006B",X"006C",X"006C",X"0068",X"0062",
    X"005F",X"0055",X"0050",X"0048",X"0042",X"0038",X"002E",X"0020",X"0018",X"000A",X"0005",X"FFF8",X"FFF0",X"FFE8",X"FFDD",X"FFD6",
    X"FFCF",X"FFCB",X"FFC8",X"FFC5",X"FFC3",X"FFC6",X"FFC8",X"FFCD",X"FFD2",X"FFD8",X"FFDF",X"FFE5",X"FFEE",X"FFF5",X"FFFF",X"0008",
    X"000E",X"0016",X"001D",X"0026",X"002D",X"0032",X"0037",X"003C",X"0040",X"0040",X"0044",X"0042",X"0043",X"0040",X"003B",X"0037",
    X"0031",X"002D",X"0023",X"001E",X"0015",X"000B",X"FFFF",X"FFF7",X"FFEC",X"FFE4",X"FFDC",X"FFD4",X"FFCD",X"FFC7",X"FFC0",X"FFBA",
    X"FFB5",X"FFB4",X"FFB2",X"FFB0",X"FFAF",X"FFB2",X"FFB6",X"FFB7",X"FFBC",X"FFC2",X"FFC7",X"FFCE",X"FFD7",X"FFDD",X"FFE5",X"FFF0",
    X"FFF8",X"0002",X"000B",X"0014",X"001B",X"0023",X"002C",X"0031",X"0039",X"003C",X"0040",X"0043",X"0046",X"0046",X"0048",X"0046",
    X"0044",X"0041",X"003D",X"0035",X"0031",X"0029",X"0021",X"001B",X"0014",X"0009",X"0003",X"FFF7",X"FFF0",X"FFE9",X"FFE1",X"FFDB",
    X"FFD4",X"FFD0",X"FFCA",X"FFC6",X"FFC3",X"FFC1",X"FFC0",X"FFBE",X"FFBD",X"FFC0",X"FFC2",X"FFC7",X"FFCB",X"FFCF",X"FFD3",X"FFDA",
    X"FFDF",X"FFE6",X"FFED",X"FFF2",X"FFF9",X"0000",X"0004",X"000A",X"0011",X"0014",X"0019",X"001E",X"0020",X"0022",X"0024",X"0024",
    X"0027",X"0027",X"0025",X"0026",X"0024",X"0021",X"001D",X"001C",X"0019",X"0015",X"0012",X"000E",X"000A",X"0005",X"0002",X"FFFE",
    X"FFF8",X"FFF5",X"FFF3",X"FFEF",X"FFEC",X"FFEA",X"FFE9",X"FFE7",X"FFE6",X"FFE6",X"FFE7",X"FFE8",X"FFE9",X"FFEB",X"FFEB",X"FFED",
    X"FFF0",X"FFF1",X"FFF4",X"FFF6",X"FFF8",X"FFFB",X"FFFE",X"0002",X"0004",X"0006",X"0008",X"0009",X"000B",X"000A",X"000A",X"000A",
    X"000B",X"000B",X"000A",X"0008",X"0007",X"0005",X"0003",X"0000",X"0000",X"FFFD",X"FFFC",X"FFF9",X"FFF7",X"FFF6",X"FFF3",X"FFF2",
    X"FFEF",X"FFEE",X"FFEC",X"FFEB",X"FFE9",X"FFE8",X"FFE9",X"FFE8",X"FFEA",X"FFEA",X"FFEA",X"FFEC",X"FFEC",X"FFEF",X"FFF1",X"FFF2",
    X"FFF4",X"FFF6",X"FFF7",X"FFF9",X"FFFA",X"FFFD",X"FFFE",X"FFFF",X"0001",X"0002",X"0004",X"0003",X"0004",X"0005",X"0007",X"0007",
    X"0007",X"0008",X"0008",X"0008",X"0007",X"0006",X"0006",X"0006",X"0004",X"0003",X"0003",X"0002",X"0001",X"FFFF",X"FFFE",X"FFFE",
    X"FFFD",X"FFFC",X"FFFC",X"FFFC",X"FFFB",X"FFFB",X"FFFB",X"FFFC",X"FFFD",X"FFFD",X"FFFF",X"0000",X"0001",X"0002",X"0002",X"0003",
    X"0004",X"0004",X"0005",X"0006",X"0008",X"0008",X"0009",X"0009",X"000B",X"000B",X"000C",X"000C",X"000C",X"000B",X"000A",X"000A",
    X"0008",X"0007",X"0006",X"0003",X"0002",X"0000",X"FFFE",X"FFFD",X"FFFA",X"FFF9",X"FFF7",X"FFF6",X"FFF5",X"FFF4",X"FFF2",X"FFF1",
    X"FFF1",X"FFF1",X"FFF0",X"FFEF",X"FFEF",X"FFF0",X"FFEF",X"FFF0",X"FFF1",X"FFF2",X"FFF4",X"FFF5",X"FFF7",X"FFF8",X"FFFA",X"FFFC",
    X"FFFD",X"FFFE",X"0000",X"0002",X"0003",X"0004",X"0006",X"0006",X"0008",X"0008",X"000A",X"000B",X"000C",X"000C",X"000D",X"000D",
    X"000D",X"000D",X"000C",X"000C",X"000B",X"000B",X"000A",X"0009",X"0008",X"0006",X"0006",X"0004",X"0002",X"0001",X"0001",X"0000",
    X"FFFF",X"FFFE",X"FFFE",X"FFFD",X"FFFD",X"FFFD",X"FFFC",X"FFFC",X"FFFC",X"FFFC",X"FFFC",X"FFFC",X"FFFD",X"FFFD",X"FFFE",X"FFFE",
    X"FFFE",X"FFFE",X"FFFF",X"0000",X"0001",X"0001",X"0002",X"0002",X"0002",X"0003",X"0004",X"0004",X"0004",X"0004",X"0005",X"0005",
    X"0004",X"0004",X"0004",X"0003",X"0003",X"0002",X"0002",X"0002",X"0002",X"0001",X"0001",X"0001",X"0000",X"FFFF",X"FFFF",X"FFFE",
    X"FFFE",X"FFFE",X"FFFD",X"FFFD",X"FFFC",X"FFFC",X"FFFD",X"FFFD",X"FFFD",X"FFFD",X"FFFD",X"FFFD",X"FFFE",X"FFFE",X"FFFF",X"0000",
    X"0000",X"0001",X"0001",X"0001",X"0002",X"0002",X"0003",X"0003",X"0003",X"0003",X"0003",X"0003",X"0003",X"0003",X"0003",X"0003",
    X"0002",X"0002",X"0002",X"0002",X"0001",X"0000",X"0000",X"0000",X"FFFF",X"FFFE",X"FFFE",X"FFFD",X"FFFC",X"FFFC",X"FFFB",X"FFFA",
    X"FFFA",X"FFFA",X"FFFA",X"FFFA",X"FFF9",X"FFF9",X"FFF9",X"FFF9",X"FFF9",X"FFFA",X"FFFA",X"FFFA",X"FFFA",X"FFFB",X"FFFC",X"FFFD",
    X"FFFD",X"FFFE",X"FFFF",X"FFFF",X"0000",X"0001",X"0002",X"0002",X"0004",X"0004",X"0005",X"0005",X"0006",X"0006",X"0007",X"0007",
    X"0007",X"0008",X"0008",X"0008",X"0007",X"0007",X"0007",X"0007",X"0006",X"0006",X"0005",X"0005",X"0004",X"0003",X"0003",X"0002",
    X"0001",X"0001",X"0000",X"FFFF",X"FFFE",X"FFFE",X"FFFD",X"FFFC",X"FFFC",X"FFFB",X"FFFA",X"FFFA",X"FFF9",X"FFF9",X"FFF9",X"FFF9",
    X"FFF9",X"FFF9",X"FFF9",X"FFF9",X"FFFA",X"FFFA",X"FFFB",X"FFFB",X"FFFB",X"FFFC",X"FFFC",X"FFFD",X"FFFD",X"FFFE",X"FFFF",X"0000"
  );
begin
  process(clock) is
  begin
    if rising_edge(clock) then
      data0_1 <= WAVEFORM_DATA(to_integer(unsigned(addr0_0)));
      data1_1 <= WAVEFORM_DATA(to_integer(unsigned(addr1_0)));
    end if;
  end process;
end waveform_data;
