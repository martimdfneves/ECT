----------------------------------------------------------------------------------------------------------------------------------------------------------------
-- LSD.TOS, April 2018 (DO NOT REMOVE THIS LINE), VHDL 2008
--
-- 16x16 font (in bold face) with 128 characters.
--
-- Source (public domain):
--   MBWK
--   http://www.rinkydinkelectronics.com/r_fonts.php
--   arial_bold.c
--
-- Modified, expanded to 128 characters, and converted to VHDL.
--
-- A simple example of the use of the font_16x16_bold entity can be found in the ???_example_tl.vhd
--

library IEEE;
use     IEEE.STD_LOGIC_1164.ALL;
use     IEEE.NUMERIC_STD.ALL;

entity font_16x16_bold is
  port
  (
    clock : in std_logic; -- main clock

    char_0   : in  std_logic_vector(6 downto 0); -- character number encoded as a std_logic_vector
    row_0    : in  std_logic_vector(3 downto 0); -- row number encoded as a std_logic_vector: 0 (top) to 15 (bottom)
    column_0 : in  std_logic_vector(3 downto 0); -- column number encoded as a std_logic_vector: 0 (left) to 15 (right)
    data_1   : out std_logic                     -- pixel color ('0' means background color, '1' means foreground color)
  );
end font_16x16_bold;

architecture font_data of font_16x16_bold is
  signal addr_0x : std_logic_vector(14 downto 0); -- equal to 256*char+16*row+col
  --
  -- Single port ROM memory data
  --
  type rom_t is array(0 to 128*16*16-1) of std_logic;
  constant FONT_DATA : rom_t :=
  -- [  0,"0000000",0x00] top-left of a table box
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000001111111111" &
    "0000001111111111" &
    "0000001111111111" &
    "0000001111111111" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
  -- [  1,"0000001",0x01] top-center of a table box
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "1111111111111111" &
    "1111111111111111" &
    "1111111111111111" &
    "1111111111111111" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
  -- [  2,"0000010",0x02] top-right of a table box
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "1111111111000000" &
    "1111111111000000" &
    "1111111111000000" &
    "1111111111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
  -- [  3,"0000011",0x03] middle-left of a table box
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111111111" &
    "0000001111111111" &
    "0000001111111111" &
    "0000001111111111" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
  -- [  4,"0000100",0x04] middle-center of a table box
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "1111111111111111" &
    "1111111111111111" &
    "1111111111111111" &
    "1111111111111111" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
  -- [  5,"0000101",0x05] middle-right of a table box
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "1111111111000000" &
    "1111111111000000" &
    "1111111111000000" &
    "1111111111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
  -- [  6,"0000110",0x06] bottom-left of a table box
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111111111" &
    "0000001111111111" &
    "0000001111111111" &
    "0000001111111111" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [  7,"0000111",0x07] bottom-center of a table box
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "1111111111111111" &
    "1111111111111111" &
    "1111111111111111" &
    "1111111111111111" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [  8,"0001000",0x08] bottom-right of a table box
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "1111111111000000" &
    "1111111111000000" &
    "1111111111000000" &
    "1111111111000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [  9,"0001001",0x09] horizontal line of a table box
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "1111111111111111" &
    "1111111111111111" &
    "1111111111111111" &
    "1111111111111111" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 10,"0001010",0x0A] vertical line of a table box
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
  -- [ 11,"0001011",0x0B] rounded top-left of a table box
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000011111111" &
    "0000000111111111" &
    "0000001111111111" &
    "0000001111111111" &
    "0000001111100000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
  -- [ 12,"0001100",0x0C] rounded top-right of a table box
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "1111111100000000" &
    "1111111110000000" &
    "1111111111000000" &
    "1111111111000000" &
    "0000011111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
  -- [ 13,"0001101",0x0D] rounded bottom-left of a table box
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111100000" &
    "0000001111111111" &
    "0000001111111111" &
    "0000000111111111" &
    "0000000011111111" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 14,"0001110",0x0E] rounded bottom-right of a table box
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000011111000000" &
    "1111111111000000" &
    "1111111111000000" &
    "1111111110000000" &
    "1111111100000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 15,"0001111",0x0F] thin X inside a box
    "1111111111111111" &
    "1100000000000011" &
    "1010000000000101" &
    "1001000000001001" &
    "1000100000010001" &
    "1000010000100001" &
    "1000001001000001" &
    "1000000110000001" &
    "1000000110000001" &
    "1000001001000001" &
    "1000010000100001" &
    "1000100000010001" &
    "1001000000001001" &
    "1010000000000101" &
    "1100000000000011" &
    "1111111111111111" &
  -- [ 16,"0010000",0x10] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 17,"0010001",0x11] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 18,"0010010",0x12] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 19,"0010011",0x13] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 20,"0010100",0x14] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 21,"0010101",0x15] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 22,"0010110",0x16] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 23,"0010111",0x17] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 24,"0011000",0x18] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 25,"0011001",0x19] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 26,"0011010",0x1A] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 27,"0011011",0x1B] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 28,"0011100",0x1C] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 29,"0011101",0x1D] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 30,"0011110",0x1E] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 31,"0011111",0x1F] unused (blank)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 32,"0100000",0x20] space
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 33,"0100001",0x21] !
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 34,"0100010",0x22] "
    "0000000000000000" &
    "0000000000000000" &
    "0000011001100000" &
    "0000011001100000" &
    "0000011001100000" &
    "0000011001100000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 35,"0100011",0x23] #
    "0000000000000000" &
    "0000000000000000" &
    "0000000110110000" &
    "0000000110110000" &
    "0000001101100000" &
    "0001111111111000" &
    "0001111111111000" &
    "0000001101100000" &
    "0000011011000000" &
    "0001111111111000" &
    "0001111111111000" &
    "0000011011000000" &
    "0000110110000000" &
    "0000110110000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 36,"0100100",0x24] $
    "0000000000000000" &
    "0000000100000000" &
    "0000001110000000" &
    "0000011111000000" &
    "0000110101100000" &
    "0000110100000000" &
    "0000111100000000" &
    "0000011110000000" &
    "0000001111000000" &
    "0000000111100000" &
    "0000110101100000" &
    "0000110101100000" &
    "0000011111000000" &
    "0000001110000000" &
    "0000000100000000" &
    "0000000000000000" &
  -- [ 37,"0100101",0x25] %
    "0000000000000000" &
    "0000000000000000" &
    "0011110000011000" &
    "0110011000110000" &
    "0110011001100000" &
    "0110011001100000" &
    "0011110011000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000001100111100" &
    "0000011001100110" &
    "0000011001100110" &
    "0000110001100110" &
    "0001100000111100" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 38,"0100110",0x26] &
    "0000000000000000" &
    "0000000000000000" &
    "0000111110000000" &
    "0001111111000000" &
    "0001100011000000" &
    "0001100011000000" &
    "0000111110000000" &
    "0000111100000000" &
    "0001101100100000" &
    "0011001110110000" &
    "0011000111100000" &
    "0011000011110000" &
    "0001111111111000" &
    "0000111100010000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 39,"0100111",0x27] '
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 40,"0101000",0x28] (
    "0000000000000000" &
    "0000000000000000" &
    "0000000011000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000011000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 41,"0101001",0x29] )
    "0000000000000000" &
    "0000000000000000" &
    "0000001100000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000011000000" &
    "0000000011000000" &
    "0000000011000000" &
    "0000000011000000" &
    "0000000011000000" &
    "0000000011000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000001100000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 42,"0101010",0x2A] *
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000001110000000" &
    "0000001110000000" &
    "0011001110011000" &
    "0011111111111000" &
    "0000011111000000" &
    "0000011111000000" &
    "0000111011100000" &
    "0001110001110000" &
    "0000010001000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 43,"0101011",0x2B] +
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000111111110000" &
    "0000111111110000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 44,"0101100",0x2C] ,
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000010000000" &
    "0000000010000000" &
    "0000000100000000" &
  -- [ 45,"0101101",0x2D] -
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000011111100000" &
    "0000011111100000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 46,"0101110",0x2E] .
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 47,"0101111",0x2F] /
    "0000000000000000" &
    "0000000000000000" &
    "0000000000011000" &
    "0000000000110000" &
    "0000000001100000" &
    "0000000001100000" &
    "0000000011000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000001100000000" &
    "0000011000000000" &
    "0000011000000000" &
    "0000110000000000" &
    "0001100000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 48,"0110000",0x30] 0
    "0000000000000000" &
    "0000000000000000" &
    "0000001111000000" &
    "0000011111100000" &
    "0000111001110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000111001110000" &
    "0000011111100000" &
    "0000001111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 49,"0110001",0x31] 1
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000001110000000" &
    "0000011110000000" &
    "0000110110000000" &
    "0000100110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 50,"0110010",0x32] 2
    "0000000000000000" &
    "0000000000000000" &
    "0000001111000000" &
    "0000011111100000" &
    "0000111000110000" &
    "0000110000110000" &
    "0000000000110000" &
    "0000000001100000" &
    "0000000011100000" &
    "0000000111000000" &
    "0000001110000000" &
    "0000011000000000" &
    "0000111111110000" &
    "0000111111110000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 51,"0110011",0x33] 3
    "0000000000000000" &
    "0000000000000000" &
    "0000001111100000" &
    "0000011111110000" &
    "0000111000110000" &
    "0000000000110000" &
    "0000000111100000" &
    "0000000111100000" &
    "0000000001110000" &
    "0000000000110000" &
    "0000110000110000" &
    "0000111001110000" &
    "0000011111100000" &
    "0000001111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 52,"0110100",0x34] 4
    "0000000000000000" &
    "0000000000000000" &
    "0000000001100000" &
    "0000000011100000" &
    "0000000011100000" &
    "0000000111100000" &
    "0000001101100000" &
    "0000001101100000" &
    "0000011001100000" &
    "0000110001100000" &
    "0000111111110000" &
    "0000111111110000" &
    "0000000001100000" &
    "0000000001100000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 53,"0110101",0x35] 5
    "0000000000000000" &
    "0000000000000000" &
    "0000011111100000" &
    "0000011111100000" &
    "0000011000000000" &
    "0000110000000000" &
    "0000111111000000" &
    "0000111111100000" &
    "0000000001110000" &
    "0000000000110000" &
    "0000110000110000" &
    "0000111001110000" &
    "0000011111100000" &
    "0000001111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 54,"0110110",0x36] 6
    "0000000000000000" &
    "0000000000000000" &
    "0000001111100000" &
    "0000011111110000" &
    "0000011000110000" &
    "0000110000000000" &
    "0000110111000000" &
    "0000111111100000" &
    "0000111001110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000011000110000" &
    "0000011111100000" &
    "0000001111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 55,"0110111",0x37] 7
    "0000000000000000" &
    "0000000000000000" &
    "0000111111110000" &
    "0000111111110000" &
    "0000000001100000" &
    "0000000011000000" &
    "0000000011000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000001110000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 56,"0111000",0x38] 8
    "0000000000000000" &
    "0000000000000000" &
    "0000001111000000" &
    "0000011111100000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000011111100000" &
    "0000011111100000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000011111100000" &
    "0000001111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 57,"0111001",0x39] 9
    "0000000000000000" &
    "0000000000000000" &
    "0000001111000000" &
    "0000011111100000" &
    "0000110001100000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000111001110000" &
    "0000011111110000" &
    "0000001110110000" &
    "0000000000110000" &
    "0000110001100000" &
    "0000111111100000" &
    "0000011111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 58,"0111010",0x3A] :
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 59,"0111011",0x3B] ;
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000010000000" &
    "0000000010000000" &
    "0000000100000000" &
  -- [ 60,"0111100",0x3C] <
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000010000" &
    "0000000001110000" &
    "0000000111100000" &
    "0000011110000000" &
    "0000111000000000" &
    "0000011110000000" &
    "0000000111100000" &
    "0000000001110000" &
    "0000000000010000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 61,"0111101",0x3D] =
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0001111111110000" &
    "0001111111110000" &
    "0000000000000000" &
    "0000000000000000" &
    "0001111111110000" &
    "0001111111110000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 62,"0111110",0x3E] >
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000100000000000" &
    "0000111000000000" &
    "0000011110000000" &
    "0000000111100000" &
    "0000000001110000" &
    "0000000111100000" &
    "0000011110000000" &
    "0000111000000000" &
    "0000100000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 63,"0111111",0x3F] ?
    "0000000000000000" &
    "0000000000000000" &
    "0000001111000000" &
    "0000011111100000" &
    "0000111000110000" &
    "0000110000110000" &
    "0000000001110000" &
    "0000000011100000" &
    "0000000111000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 64,"1000000",0x40] @
    "0000000000000000" &
    "0000000000000000" &
    "0000011111000000" &
    "0000110000110000" &
    "0001001101111000" &
    "0001011111101000" &
    "0010110011001000" &
    "0010110011001000" &
    "0010110011001000" &
    "0010111111010000" &
    "0010011011100000" &
    "0001000000001000" &
    "0000100000010000" &
    "0000011111100000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 65,"1000001",0x41] A
    "0000000000000000" &
    "0000000000000000" &
    "0000001110000000" &
    "0000001110000000" &
    "0000011011000000" &
    "0000011011000000" &
    "0000011011000000" &
    "0000110001100000" &
    "0000110001100000" &
    "0000111111100000" &
    "0001111111110000" &
    "0001100000110000" &
    "0001100000110000" &
    "0011000000011000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 66,"1000010",0x42] B
    "0000000000000000" &
    "0000000000000000" &
    "0001111111100000" &
    "0001111111110000" &
    "0001100000110000" &
    "0001100000110000" &
    "0001100000110000" &
    "0001111111100000" &
    "0001111111110000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001111111110000" &
    "0001111111100000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 67,"1000011",0x43] C
    "0000000000000000" &
    "0000000000000000" &
    "0000001111100000" &
    "0000111111110000" &
    "0000110000111000" &
    "0001110000010000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001110000010000" &
    "0000110000111000" &
    "0000111111110000" &
    "0000001111100000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 68,"1000100",0x44] D
    "0000000000000000" &
    "0000000000000000" &
    "0001111111000000" &
    "0001111111110000" &
    "0001100000110000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000110000" &
    "0001111111110000" &
    "0001111111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 69,"1000101",0x45] E
    "0000000000000000" &
    "0000000000000000" &
    "0001111111111000" &
    "0001111111111000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001111111111000" &
    "0001111111111000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001111111111000" &
    "0001111111111000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 70,"1000110",0x46] F
    "0000000000000000" &
    "0000000000000000" &
    "0001111111111000" &
    "0001111111111000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001111111000000" &
    "0001111111000000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001100000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 71,"1000111",0x47] G
    "0000000000000000" &
    "0000000000000000" &
    "0000011111100000" &
    "0001111111110000" &
    "0001100000111000" &
    "0011100000010000" &
    "0011000000000000" &
    "0011000000000000" &
    "0011000011111000" &
    "0011000011111000" &
    "0011100000011000" &
    "0001100000111000" &
    "0001111111111000" &
    "0000011111100000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 72,"1001000",0x48] H
    "0000000000000000" &
    "0000000000000000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001111111111000" &
    "0001111111111000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 73,"1001001",0x49] I
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 74,"1001010",0x4A] J
    "0000000000000000" &
    "0000000000000000" &
    "0000000000110000" &
    "0000000000110000" &
    "0000000000110000" &
    "0000000000110000" &
    "0000000000110000" &
    "0000000000110000" &
    "0000000000110000" &
    "0000000000110000" &
    "0000110000110000" &
    "0000111001110000" &
    "0000011111100000" &
    "0000001111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 75,"1001011",0x4B] K
    "0000000000000000" &
    "0000000000000000" &
    "0001100000011000" &
    "0001100000110000" &
    "0001100001100000" &
    "0001100011000000" &
    "0001100110000000" &
    "0001101111000000" &
    "0001111011000000" &
    "0001110001100000" &
    "0001100001110000" &
    "0001100000110000" &
    "0001100000011000" &
    "0001100000011000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 76,"1001100",0x4C] L
    "0000000000000000" &
    "0000000000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000111111110000" &
    "0000111111110000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 77,"1001101",0x4D] M
    "0000000000000000" &
    "0000000000000000" &
    "0011100000111000" &
    "0011100000111000" &
    "0011110001111000" &
    "0011110001111000" &
    "0011010001011000" &
    "0011011011011000" &
    "0011011011011000" &
    "0011011011011000" &
    "0011001110011000" &
    "0011001110011000" &
    "0011001110011000" &
    "0011000100011000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 78,"1001110",0x4E] N
    "0000000000000000" &
    "0000000000000000" &
    "0001100000011000" &
    "0001110000011000" &
    "0001111000011000" &
    "0001111000011000" &
    "0001101100011000" &
    "0001100110011000" &
    "0001100110011000" &
    "0001100011011000" &
    "0001100001111000" &
    "0001100001111000" &
    "0001100000111000" &
    "0001100000011000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 79,"1001111",0x4F] O
    "0000000000000000" &
    "0000000000000000" &
    "0000011111000000" &
    "0001111111110000" &
    "0001100000110000" &
    "0011000000011000" &
    "0011000000011000" &
    "0011000000011000" &
    "0011000000011000" &
    "0011000000011000" &
    "0011000000011000" &
    "0001100000110000" &
    "0001111111110000" &
    "0000011111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 80,"1010000",0x50] P
    "0000000000000000" &
    "0000000000000000" &
    "0001111111000000" &
    "0001111111100000" &
    "0001100001110000" &
    "0001100000110000" &
    "0001100001110000" &
    "0001111111100000" &
    "0001111111000000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001100000000000" &
    "0001100000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 81,"1010001",0x51] Q
    "0000000000000000" &
    "0000000000000000" &
    "0000011111000000" &
    "0001111111110000" &
    "0001100000110000" &
    "0011000000011000" &
    "0011000000011000" &
    "0011000000011000" &
    "0011000000011000" &
    "0011000000011000" &
    "0011000110111000" &
    "0001100011110000" &
    "0001111111110000" &
    "0000011110110000" &
    "0000000000011000" &
    "0000000000000000" &
  -- [ 82,"1010010",0x52] R
    "0000000000000000" &
    "0000000000000000" &
    "0001111111100000" &
    "0001111111110000" &
    "0001100000111000" &
    "0001100000011000" &
    "0001100000111000" &
    "0001111111110000" &
    "0001111111000000" &
    "0001100011100000" &
    "0001100001110000" &
    "0001100000110000" &
    "0001100000111000" &
    "0001100000011100" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 83,"1010011",0x53] S
    "0000000000000000" &
    "0000000000000000" &
    "0000011111000000" &
    "0000111111100000" &
    "0001110001110000" &
    "0001100000110000" &
    "0001111000000000" &
    "0000111111000000" &
    "0000001111100000" &
    "0000000001110000" &
    "0001100000110000" &
    "0001110001110000" &
    "0000111111100000" &
    "0000011111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 84,"1010100",0x54] T
    "0000000000000000" &
    "0000000000000000" &
    "0001111111111000" &
    "0001111111111000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 85,"1010101",0x55] U
    "0000000000000000" &
    "0000000000000000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001100000011000" &
    "0001110000111000" &
    "0000111111110000" &
    "0000011111100000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 86,"1010110",0x56] V
    "0000000000000000" &
    "0000000000000000" &
    "0011000000011000" &
    "0001100000110000" &
    "0001100000110000" &
    "0001100000110000" &
    "0000110001100000" &
    "0000110001100000" &
    "0000111011100000" &
    "0000011011000000" &
    "0000011011000000" &
    "0000001110000000" &
    "0000001110000000" &
    "0000001110000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 87,"1010111",0x57] W
    "0000000000000000" &
    "0000000000000000" &
    "0011000111000110" &
    "0011000111000110" &
    "0011000111000110" &
    "0001101101101100" &
    "0001101101101100" &
    "0001101101101100" &
    "0001101101101100" &
    "0001101101101100" &
    "0000111000111000" &
    "0000111000111000" &
    "0000111000111000" &
    "0000111000111000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 88,"1011000",0x58] X
    "0000000000000000" &
    "0000000000000000" &
    "0001100000110000" &
    "0001110001110000" &
    "0000110001100000" &
    "0000011011000000" &
    "0000011111000000" &
    "0000001110000000" &
    "0000001110000000" &
    "0000011111000000" &
    "0000011011000000" &
    "0000110001100000" &
    "0001110001110000" &
    "0001100000110000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 89,"1011001",0x59] Y
    "0000000000000000" &
    "0000000000000000" &
    "0001100000011000" &
    "0001110000111000" &
    "0000110000110000" &
    "0000011001100000" &
    "0000011001100000" &
    "0000001111000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 90,"1011010",0x5A] Z
    "0000000000000000" &
    "0000000000000000" &
    "0000111111110000" &
    "0000111111110000" &
    "0000000001100000" &
    "0000000011000000" &
    "0000000111000000" &
    "0000000110000000" &
    "0000001100000000" &
    "0000011100000000" &
    "0000011000000000" &
    "0000110000000000" &
    "0001111111110000" &
    "0001111111110000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 91,"1011011",0x5B] [
    "0000000000000000" &
    "0000000000000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 92,"1011100",0x5C] \
    "0000000000000000" &
    "0000000000000000" &
    "0001100000000000" &
    "0000110000000000" &
    "0000011000000000" &
    "0000011000000000" &
    "0000001100000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000011000000" &
    "0000000001100000" &
    "0000000001100000" &
    "0000000000110000" &
    "0000000000011000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 93,"1011101",0x5D] ]
    "0000000000000000" &
    "0000000000000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000000011000000" &
    "0000000011000000" &
    "0000000011000000" &
    "0000000011000000" &
    "0000000011000000" &
    "0000000011000000" &
    "0000000011000000" &
    "0000000011000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 94,"1011110",0x5E] ^
    "0000000000000000" &
    "0000000110000000" &
    "0000001111000000" &
    "0000001111000000" &
    "0000011001100000" &
    "0000011001100000" &
    "0000011001100000" &
    "0000110000110000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 95,"1011111",0x5F] _
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0011111111111100" &
    "0011111111111100" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 96,"1100000",0x60] `
    "0000000000000000" &
    "0000000000000000" &
    "0000001100000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 97,"1100001",0x61] a
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000011111000000" &
    "0000111111100000" &
    "0000110001100000" &
    "0000000111100000" &
    "0000011111100000" &
    "0000111001100000" &
    "0000110001100000" &
    "0000111111100000" &
    "0000011110110000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 98,"1100010",0x62] b
    "0000000000000000" &
    "0000000000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110111000000" &
    "0000111111100000" &
    "0000111001110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000111001110000" &
    "0000111111100000" &
    "0000110111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [ 99,"1100011",0x63] c
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000001111000000" &
    "0000011111100000" &
    "0000111001100000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000111001100000" &
    "0000011111100000" &
    "0000001111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [100,"1100100",0x64] d
    "0000000000000000" &
    "0000000000000000" &
    "0000000000110000" &
    "0000000000110000" &
    "0000000000110000" &
    "0000001110110000" &
    "0000011111110000" &
    "0000111001110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000111001110000" &
    "0000011111110000" &
    "0000001110110000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [101,"1100101",0x65] e
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000001110000000" &
    "0000011111000000" &
    "0000110001100000" &
    "0000111111100000" &
    "0000111111100000" &
    "0000110000000000" &
    "0000111001100000" &
    "0000011111000000" &
    "0000001110000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [102,"1100110",0x66] f
    "0000000000000000" &
    "0000000000000000" &
    "0000001111000000" &
    "0000011111000000" &
    "0000011000000000" &
    "0000111110000000" &
    "0000111110000000" &
    "0000011000000000" &
    "0000011000000000" &
    "0000011000000000" &
    "0000011000000000" &
    "0000011000000000" &
    "0000011000000000" &
    "0000011000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [103,"1100111",0x67] g
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000011101100000" &
    "0000111111100000" &
    "0001110011100000" &
    "0001100001100000" &
    "0001100001100000" &
    "0001100001100000" &
    "0001110011100000" &
    "0000111111100000" &
    "0000011101100000" &
    "0001100001100000" &
    "0001111111100000" &
    "0000111111000000" &
  -- [104,"1101000",0x68] h
    "0000000000000000" &
    "0000000000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110111100000" &
    "0000111111110000" &
    "0000111000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [105,"1101001",0x69] i
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [106,"1101010",0x6A] j
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000011110000000" &
    "0000011100000000" &
  -- [107,"1101011",0x6B] k
    "0000000000000000" &
    "0000000000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110000000000" &
    "0000110001100000" &
    "0000110011000000" &
    "0000110110000000" &
    "0000111110000000" &
    "0000111111000000" &
    "0000111011000000" &
    "0000110011000000" &
    "0000110001100000" &
    "0000110001100000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [108,"1101100",0x6C] l
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000011000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [109,"1101101",0x6D] m
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0011011100111000" &
    "0011111111111100" &
    "0011100111001100" &
    "0011000110001100" &
    "0011000110001100" &
    "0011000110001100" &
    "0011000110001100" &
    "0011000110001100" &
    "0011000110001100" &
    "0000000000000000" &
    "0000000000000000" &
  -- [110,"1101110",0x6E] n
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000110111100000" &
    "0000111111110000" &
    "0000111000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [111,"1101111",0x6F] o
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000001111000000" &
    "0000011111100000" &
    "0000111001110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000111001110000" &
    "0000011111100000" &
    "0000001111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [112,"1110000",0x70] p
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000110111000000" &
    "0000111111100000" &
    "0000111001110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000111001110000" &
    "0000111111100000" &
    "0000110111000000" &
    "0000110000000000" &
    "0000110000000000" &
  -- [113,"1110001",0x71] q
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000001110110000" &
    "0000011111110000" &
    "0000111001110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000111001110000" &
    "0000011111110000" &
    "0000001110110000" &
    "0000000000110000" &
    "0000000000110000" &
  -- [114,"1110010",0x72] r
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000001101110000" &
    "0000001111110000" &
    "0000001110000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [115,"1110011",0x73] s
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000011111000000" &
    "0000111111100000" &
    "0000110001100000" &
    "0000111100000000" &
    "0000011111000000" &
    "0000000011100000" &
    "0000110001100000" &
    "0000111111100000" &
    "0000011111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [116,"1110100",0x74] t
    "0000000000000000" &
    "0000000000000000" &
    "0000000100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000011111000000" &
    "0000011111000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001100000000" &
    "0000001111000000" &
    "0000000111000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [117,"1110101",0x75] u
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110000110000" &
    "0000110001110000" &
    "0000111111110000" &
    "0000011110110000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [118,"1110110",0x76] v
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000110001100000" &
    "0000110001100000" &
    "0000110001100000" &
    "0000011011000000" &
    "0000011011000000" &
    "0000011011000000" &
    "0000001110000000" &
    "0000001110000000" &
    "0000001110000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [119,"1110111",0x77] w
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0011000111000110" &
    "0011000111000110" &
    "0001100111001100" &
    "0001101101101100" &
    "0001101101101100" &
    "0001101101101100" &
    "0000111000111000" &
    "0000111000111000" &
    "0000111000111000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [120,"1111000",0x78] x
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000011000110000" &
    "0000011101110000" &
    "0000001101100000" &
    "0000000111000000" &
    "0000000111000000" &
    "0000000111000000" &
    "0000001101100000" &
    "0000011101110000" &
    "0000011000110000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [121,"1111001",0x79] y
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000110000011000" &
    "0000110000011000" &
    "0000011000110000" &
    "0000011000110000" &
    "0000001101100000" &
    "0000001101100000" &
    "0000001111100000" &
    "0000000111000000" &
    "0000000111000000" &
    "0000000110000000" &
    "0000011110000000" &
    "0000011100000000" &
  -- [122,"1111010",0x7A] z
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000111111100000" &
    "0000111111100000" &
    "0000000011000000" &
    "0000000111000000" &
    "0000001110000000" &
    "0000011100000000" &
    "0000011000000000" &
    "0000111111100000" &
    "0000111111100000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [123,"1111011",0x7B] {
    "0000000000000000" &
    "0000000000000000" &
    "0000000011100000" &
    "0000000111100000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000011100000000" &
    "0000011100000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000111100000" &
    "0000000011100000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [124,"1111100",0x7C] |
    "0000000000000000" &
    "0000000000000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [125,"1111101",0x7D] }
    "0000000000000000" &
    "0000000000000000" &
    "0000011100000000" &
    "0000011110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000011100000" &
    "0000000011100000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000000110000000" &
    "0000011110000000" &
    "0000011100000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [126,"1111110",0x7E] ~
    "0000000000000000" &
    "0000000000000000" &
    "0000111100010000" &
    "0001111111110000" &
    "0001000111100000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
  -- [127,"1111111",0x7F] filled o (a disk)
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000000000000000" &
    "0000001111000000" &
    "0000011111100000" &
    "0000111111110000" &
    "0000111111110000" &
    "0000111111110000" &
    "0000111111110000" &
    "0000111111110000" &
    "0000011111100000" &
    "0000001111000000" &
    "0000000000000000" &
    "0000000000000000";
begin
  addr_0x <= char_0 & row_0 & column_0;
  process(clock) is
  begin
    if rising_edge(clock) then
      data_1 <= FONT_DATA(to_integer(unsigned(addr_0x)));
    end if;
  end process;
end font_data;
